// int32 mul
// deyuan, 09/25/2024

module mul_int32(input [3:0] pi0, input [3:0] pi1, output [3:0] po0);
    assign po0 = pi0 * pi1;
endmodule

