// AES sbox
// hosein, 09/17/2024

module sbox(input [7:0] pi0, output reg[7:0] po0);

always @(*) begin
    case( pi0 )

        8'h00: po0 = 8'h63;
		8'h01: po0 = 8'h7C;
		8'h02: po0 = 8'h77;
		8'h03: po0 = 8'h7B;
		8'h04: po0 = 8'hF2;
		8'h05: po0 = 8'h6B;
		8'h06: po0 = 8'h6F;
		8'h07: po0 = 8'hC5;
		8'h08: po0 = 8'h30;
		8'h09: po0 = 8'h01;
		8'h0A: po0 = 8'h67;
		8'h0B: po0 = 8'h2B;
		8'h0C: po0 = 8'hFE;
		8'h0D: po0 = 8'hD7;
		8'h0E: po0 = 8'hAB;
		8'h0F: po0 = 8'h76;
		8'h10: po0 = 8'hCA;
		8'h11: po0 = 8'h82;
		8'h12: po0 = 8'hC9;
		8'h13: po0 = 8'h7D;
		8'h14: po0 = 8'hFA;
		8'h15: po0 = 8'h59;
		8'h16: po0 = 8'h47;
		8'h17: po0 = 8'hF0;
		8'h18: po0 = 8'hAD;
		8'h19: po0 = 8'hD4;
		8'h1A: po0 = 8'hA2;
		8'h1B: po0 = 8'hAF;
		8'h1C: po0 = 8'h9C;
		8'h1D: po0 = 8'hA4;
		8'h1E: po0 = 8'h72;
		8'h1F: po0 = 8'hC0;
		8'h20: po0 = 8'hB7;
		8'h21: po0 = 8'hFD;
		8'h22: po0 = 8'h93;
		8'h23: po0 = 8'h26;
		8'h24: po0 = 8'h36;
		8'h25: po0 = 8'h3F;
		8'h26: po0 = 8'hF7;
		8'h27: po0 = 8'hCC;
		8'h28: po0 = 8'h34;
		8'h29: po0 = 8'hA5;
		8'h2A: po0 = 8'hE5;
		8'h2B: po0 = 8'hF1;
		8'h2C: po0 = 8'h71;
		8'h2D: po0 = 8'hD8;
		8'h2E: po0 = 8'h31;
		8'h2F: po0 = 8'h15;
		8'h30: po0 = 8'h04;
		8'h31: po0 = 8'hC7;
		8'h32: po0 = 8'h23;
		8'h33: po0 = 8'hC3;
		8'h34: po0 = 8'h18;
		8'h35: po0 = 8'h96;
		8'h36: po0 = 8'h05;
		8'h37: po0 = 8'h9A;
		8'h38: po0 = 8'h07;
		8'h39: po0 = 8'h12;
		8'h3A: po0 = 8'h80;
		8'h3B: po0 = 8'hE2;
		8'h3C: po0 = 8'hEB;
		8'h3D: po0 = 8'h27;
		8'h3E: po0 = 8'hB2;
		8'h3F: po0 = 8'h75;
		8'h40: po0 = 8'h09;
		8'h41: po0 = 8'h83;
		8'h42: po0 = 8'h2C;
		8'h43: po0 = 8'h1A;
		8'h44: po0 = 8'h1B;
		8'h45: po0 = 8'h6E;
		8'h46: po0 = 8'h5A;
		8'h47: po0 = 8'hA0;
		8'h48: po0 = 8'h52;
		8'h49: po0 = 8'h3B;
		8'h4A: po0 = 8'hD6;
		8'h4B: po0 = 8'hB3;
		8'h4C: po0 = 8'h29;
		8'h4D: po0 = 8'hE3;
		8'h4E: po0 = 8'h2F;
		8'h4F: po0 = 8'h84;
		8'h50: po0 = 8'h53;
		8'h51: po0 = 8'hD1;
		8'h52: po0 = 8'h00;
		8'h53: po0 = 8'hED;
		8'h54: po0 = 8'h20;
		8'h55: po0 = 8'hFC;
		8'h56: po0 = 8'hB1;
		8'h57: po0 = 8'h5B;
		8'h58: po0 = 8'h6A;
		8'h59: po0 = 8'hCB;
		8'h5A: po0 = 8'hBE;
		8'h5B: po0 = 8'h39;
		8'h5C: po0 = 8'h4A;
		8'h5D: po0 = 8'h4C;
		8'h5E: po0 = 8'h58;
		8'h5F: po0 = 8'hCF;
		8'h60: po0 = 8'hD0;
		8'h61: po0 = 8'hEF;
		8'h62: po0 = 8'hAA;
		8'h63: po0 = 8'hFB;
		8'h64: po0 = 8'h43;
		8'h65: po0 = 8'h4D;
		8'h66: po0 = 8'h33;
		8'h67: po0 = 8'h85;
		8'h68: po0 = 8'h45;
		8'h69: po0 = 8'hF9;
		8'h6A: po0 = 8'h02;
		8'h6B: po0 = 8'h7F;
		8'h6C: po0 = 8'h50;
		8'h6D: po0 = 8'h3C;
		8'h6E: po0 = 8'h9F;
		8'h6F: po0 = 8'hA8;
		8'h70: po0 = 8'h51;
		8'h71: po0 = 8'hA3;
		8'h72: po0 = 8'h40;
		8'h73: po0 = 8'h8F;
		8'h74: po0 = 8'h92;
		8'h75: po0 = 8'h9D;
		8'h76: po0 = 8'h38;
		8'h77: po0 = 8'hF5;
		8'h78: po0 = 8'hBC;
		8'h79: po0 = 8'hB6;
		8'h7A: po0 = 8'hDA;
		8'h7B: po0 = 8'h21;
		8'h7C: po0 = 8'h10;
		8'h7D: po0 = 8'hFF;
		8'h7E: po0 = 8'hF3;
		8'h7F: po0 = 8'hD2;
		8'h80: po0 = 8'hCD;
		8'h81: po0 = 8'h0C;
		8'h82: po0 = 8'h13;
		8'h83: po0 = 8'hEC;
		8'h84: po0 = 8'h5F;
		8'h85: po0 = 8'h97;
		8'h86: po0 = 8'h44;
		8'h87: po0 = 8'h17;
		8'h88: po0 = 8'hC4;
		8'h89: po0 = 8'hA7;
		8'h8A: po0 = 8'h7E;
		8'h8B: po0 = 8'h3D;
		8'h8C: po0 = 8'h64;
		8'h8D: po0 = 8'h5D;
		8'h8E: po0 = 8'h19;
		8'h8F: po0 = 8'h73;
		8'h90: po0 = 8'h60;
		8'h91: po0 = 8'h81;
		8'h92: po0 = 8'h4F;
		8'h93: po0 = 8'hDC;
		8'h94: po0 = 8'h22;
		8'h95: po0 = 8'h2A;
		8'h96: po0 = 8'h90;
		8'h97: po0 = 8'h88;
		8'h98: po0 = 8'h46;
		8'h99: po0 = 8'hEE;
		8'h9A: po0 = 8'hB8;
		8'h9B: po0 = 8'h14;
		8'h9C: po0 = 8'hDE;
		8'h9D: po0 = 8'h5E;
		8'h9E: po0 = 8'h0B;
		8'h9F: po0 = 8'hDB;
		8'hA0: po0 = 8'hE0;
		8'hA1: po0 = 8'h32;
		8'hA2: po0 = 8'h3A;
		8'hA3: po0 = 8'h0A;
		8'hA4: po0 = 8'h49;
		8'hA5: po0 = 8'h06;
		8'hA6: po0 = 8'h24;
		8'hA7: po0 = 8'h5C;
		8'hA8: po0 = 8'hC2;
		8'hA9: po0 = 8'hD3;
		8'hAA: po0 = 8'hAC;
		8'hAB: po0 = 8'h62;
		8'hAC: po0 = 8'h91;
		8'hAD: po0 = 8'h95;
		8'hAE: po0 = 8'hE4;
		8'hAF: po0 = 8'h79;
		8'hB0: po0 = 8'hE7;
		8'hB1: po0 = 8'hC8;
		8'hB2: po0 = 8'h37;
		8'hB3: po0 = 8'h6D;
		8'hB4: po0 = 8'h8D;
		8'hB5: po0 = 8'hD5;
		8'hB6: po0 = 8'h4E;
		8'hB7: po0 = 8'hA9;
		8'hB8: po0 = 8'h6C;
		8'hB9: po0 = 8'h56;
		8'hBA: po0 = 8'hF4;
		8'hBB: po0 = 8'hEA;
		8'hBC: po0 = 8'h65;
		8'hBD: po0 = 8'h7A;
		8'hBE: po0 = 8'hAE;
		8'hBF: po0 = 8'h08;
		8'hC0: po0 = 8'hBA;
		8'hC1: po0 = 8'h78;
		8'hC2: po0 = 8'h25;
		8'hC3: po0 = 8'h2E;
		8'hC4: po0 = 8'h1C;
		8'hC5: po0 = 8'hA6;
		8'hC6: po0 = 8'hB4;
		8'hC7: po0 = 8'hC6;
		8'hC8: po0 = 8'hE8;
		8'hC9: po0 = 8'hDD;
		8'hCA: po0 = 8'h74;
		8'hCB: po0 = 8'h1F;
		8'hCC: po0 = 8'h4B;
		8'hCD: po0 = 8'hBD;
		8'hCE: po0 = 8'h8B;
		8'hCF: po0 = 8'h8A;
		8'hD0: po0 = 8'h70;
		8'hD1: po0 = 8'h3E;
		8'hD2: po0 = 8'hB5;
		8'hD3: po0 = 8'h66;
		8'hD4: po0 = 8'h48;
		8'hD5: po0 = 8'h03;
		8'hD6: po0 = 8'hF6;
		8'hD7: po0 = 8'h0E;
		8'hD8: po0 = 8'h61;
		8'hD9: po0 = 8'h35;
		8'hDA: po0 = 8'h57;
		8'hDB: po0 = 8'hB9;
		8'hDC: po0 = 8'h86;
		8'hDD: po0 = 8'hC1;
		8'hDE: po0 = 8'h1D;
		8'hDF: po0 = 8'h9E;
		8'hE0: po0 = 8'hE1;
		8'hE1: po0 = 8'hF8;
		8'hE2: po0 = 8'h98;
		8'hE3: po0 = 8'h11;
		8'hE4: po0 = 8'h69;
		8'hE5: po0 = 8'hD9;
		8'hE6: po0 = 8'h8E;
		8'hE7: po0 = 8'h94;
		8'hE8: po0 = 8'h9B;
		8'hE9: po0 = 8'h1E;
		8'hEA: po0 = 8'h87;
		8'hEB: po0 = 8'hE9;
		8'hEC: po0 = 8'hCE;
		8'hED: po0 = 8'h55;
		8'hEE: po0 = 8'h28;
		8'hEF: po0 = 8'hDF;
		8'hF0: po0 = 8'h8C;
		8'hF1: po0 = 8'hA1;
		8'hF2: po0 = 8'h89;
		8'hF3: po0 = 8'h0D;
		8'hF4: po0 = 8'hBF;
		8'hF5: po0 = 8'hE6;
		8'hF6: po0 = 8'h42;
		8'hF7: po0 = 8'h68;
		8'hF8: po0 = 8'h41;
		8'hF9: po0 = 8'h99;
		8'hFA: po0 = 8'h2D;
		8'hFB: po0 = 8'h0F;
		8'hFC: po0 = 8'hB0;
		8'hFD: po0 = 8'h54;
		8'hFE: po0 = 8'hBB;
		8'hFF: po0 = 8'h16;
        default: po0 = 0;
    endcase
end
endmodule
