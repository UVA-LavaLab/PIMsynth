// int32 div
// deyuan, 09/25/2024

module div_int32(input [31:0] a, input [31:0] b, output [31:0] q);
    assign q = a / b;
endmodule

