// int32 add
// deyuan, 09/25/2024

module add_int32(input [31:0] a, input [31:0] b, output [31:0] result);
    //assign result = a + b;
    wire n386, n387, n389, n390, n391, n392, n393, n394, n396, n397, n398,
      n399, n400, n401, n402, n404, n405, n406, n407, n408, n409, n410, n412,
      n413, n414, n415, n416, n417, n418, n420, n421, n422, n423, n424, n425,
      n426, n428, n429, n430, n431, n432, n433, n434, n436, n437, n438, n439,
      n440, n441, n442, n444, n445, n446, n447, n448, n449, n450, n452, n453,
      n454, n455, n456, n457, n458, n460, n461, n462, n463, n464, n465, n466,
      n468, n469, n470, n471, n472, n473, n474, n476, n477, n478, n479, n480,
      n481, n482, n484, n485, n486, n487, n488, n489, n490, n492, n493, n494,
      n495, n496, n497, n498, n500, n501, n502, n503, n504, n505, n506, n508,
      n509, n510, n511, n512, n513, n514, n516, n517, n518, n519, n520, n521,
      n522, n524, n525, n526, n527, n528, n529, n530, n532, n533, n534, n535,
      n536, n537, n538, n540, n541, n542, n543, n544, n545, n546, n548, n549,
      n550, n551, n552, n553, n554, n556, n557, n558, n559, n560, n561, n562,
      n564, n565, n566, n567, n568, n569, n570, n572, n573, n574, n575, n576,
      n577, n578, n580, n581, n582, n583, n584, n585, n586, n588, n589, n590,
      n591, n592, n593, n594, n596, n597, n598, n599, n600, n601, n602, n604,
      n605, n606, n607, n608, n609, n610, n612, n613, n614, n615, n616, n617,
      n618, n620, n621, n622, n623, n624, n625, n626, n628, n629, n630, n631,
      n632, n633, n634;
    assign n386 = a[0]  & ~b[0] ;
    assign n387 = ~a[0]  & b[0] ;
    assign result[0]  = n386 | n387;
    assign n389 = a[0]  & b[0] ;
    assign n390 = ~a[1]  & ~b[1] ;
    assign n391 = a[1]  & b[1] ;
    assign n392 = ~n390 & ~n391;
    assign n393 = n389 & ~n392;
    assign n394 = ~n389 & n392;
    assign result[1]  = n393 | n394;
    assign n396 = n389 & ~n390;
    assign n397 = ~n391 & ~n396;
    assign n398 = ~a[2]  & ~b[2] ;
    assign n399 = a[2]  & b[2] ;
    assign n400 = ~n398 & ~n399;
    assign n401 = n397 & ~n400;
    assign n402 = ~n397 & n400;
    assign result[2]  = ~n401 & ~n402;
    assign n404 = ~n397 & ~n398;
    assign n405 = ~n399 & ~n404;
    assign n406 = ~a[3]  & ~b[3] ;
    assign n407 = a[3]  & b[3] ;
    assign n408 = ~n406 & ~n407;
    assign n409 = n405 & ~n408;
    assign n410 = ~n405 & n408;
    assign result[3]  = ~n409 & ~n410;
    assign n412 = ~n405 & ~n406;
    assign n413 = ~n407 & ~n412;
    assign n414 = ~a[4]  & ~b[4] ;
    assign n415 = a[4]  & b[4] ;
    assign n416 = ~n414 & ~n415;
    assign n417 = n413 & ~n416;
    assign n418 = ~n413 & n416;
    assign result[4]  = ~n417 & ~n418;
    assign n420 = ~n413 & ~n414;
    assign n421 = ~n415 & ~n420;
    assign n422 = ~a[5]  & ~b[5] ;
    assign n423 = a[5]  & b[5] ;
    assign n424 = ~n422 & ~n423;
    assign n425 = n421 & ~n424;
    assign n426 = ~n421 & n424;
    assign result[5]  = ~n425 & ~n426;
    assign n428 = ~n421 & ~n422;
    assign n429 = ~n423 & ~n428;
    assign n430 = ~a[6]  & ~b[6] ;
    assign n431 = a[6]  & b[6] ;
    assign n432 = ~n430 & ~n431;
    assign n433 = n429 & ~n432;
    assign n434 = ~n429 & n432;
    assign result[6]  = ~n433 & ~n434;
    assign n436 = ~n429 & ~n430;
    assign n437 = ~n431 & ~n436;
    assign n438 = ~a[7]  & ~b[7] ;
    assign n439 = a[7]  & b[7] ;
    assign n440 = ~n438 & ~n439;
    assign n441 = n437 & ~n440;
    assign n442 = ~n437 & n440;
    assign result[7]  = ~n441 & ~n442;
    assign n444 = ~n437 & ~n438;
    assign n445 = ~n439 & ~n444;
    assign n446 = ~a[8]  & ~b[8] ;
    assign n447 = a[8]  & b[8] ;
    assign n448 = ~n446 & ~n447;
    assign n449 = n445 & ~n448;
    assign n450 = ~n445 & n448;
    assign result[8]  = ~n449 & ~n450;
    assign n452 = ~n445 & ~n446;
    assign n453 = ~n447 & ~n452;
    assign n454 = ~a[9]  & ~b[9] ;
    assign n455 = a[9]  & b[9] ;
    assign n456 = ~n454 & ~n455;
    assign n457 = n453 & ~n456;
    assign n458 = ~n453 & n456;
    assign result[9]  = ~n457 & ~n458;
    assign n460 = ~n453 & ~n454;
    assign n461 = ~n455 & ~n460;
    assign n462 = ~a[10]  & ~b[10] ;
    assign n463 = a[10]  & b[10] ;
    assign n464 = ~n462 & ~n463;
    assign n465 = n461 & ~n464;
    assign n466 = ~n461 & n464;
    assign result[10]  = ~n465 & ~n466;
    assign n468 = ~n461 & ~n462;
    assign n469 = ~n463 & ~n468;
    assign n470 = ~a[11]  & ~b[11] ;
    assign n471 = a[11]  & b[11] ;
    assign n472 = ~n470 & ~n471;
    assign n473 = n469 & ~n472;
    assign n474 = ~n469 & n472;
    assign result[11]  = ~n473 & ~n474;
    assign n476 = ~n469 & ~n470;
    assign n477 = ~n471 & ~n476;
    assign n478 = ~a[12]  & ~b[12] ;
    assign n479 = a[12]  & b[12] ;
    assign n480 = ~n478 & ~n479;
    assign n481 = n477 & ~n480;
    assign n482 = ~n477 & n480;
    assign result[12]  = ~n481 & ~n482;
    assign n484 = ~n477 & ~n478;
    assign n485 = ~n479 & ~n484;
    assign n486 = ~a[13]  & ~b[13] ;
    assign n487 = a[13]  & b[13] ;
    assign n488 = ~n486 & ~n487;
    assign n489 = n485 & ~n488;
    assign n490 = ~n485 & n488;
    assign result[13]  = ~n489 & ~n490;
    assign n492 = ~n485 & ~n486;
    assign n493 = ~n487 & ~n492;
    assign n494 = ~a[14]  & ~b[14] ;
    assign n495 = a[14]  & b[14] ;
    assign n496 = ~n494 & ~n495;
    assign n497 = n493 & ~n496;
    assign n498 = ~n493 & n496;
    assign result[14]  = ~n497 & ~n498;
    assign n500 = ~n493 & ~n494;
    assign n501 = ~n495 & ~n500;
    assign n502 = ~a[15]  & ~b[15] ;
    assign n503 = a[15]  & b[15] ;
    assign n504 = ~n502 & ~n503;
    assign n505 = n501 & ~n504;
    assign n506 = ~n501 & n504;
    assign result[15]  = ~n505 & ~n506;
    assign n508 = ~n501 & ~n502;
    assign n509 = ~n503 & ~n508;
    assign n510 = ~a[16]  & ~b[16] ;
    assign n511 = a[16]  & b[16] ;
    assign n512 = ~n510 & ~n511;
    assign n513 = n509 & ~n512;
    assign n514 = ~n509 & n512;
    assign result[16]  = ~n513 & ~n514;
    assign n516 = ~n509 & ~n510;
    assign n517 = ~n511 & ~n516;
    assign n518 = ~a[17]  & ~b[17] ;
    assign n519 = a[17]  & b[17] ;
    assign n520 = ~n518 & ~n519;
    assign n521 = n517 & ~n520;
    assign n522 = ~n517 & n520;
    assign result[17]  = ~n521 & ~n522;
    assign n524 = ~n517 & ~n518;
    assign n525 = ~n519 & ~n524;
    assign n526 = ~a[18]  & ~b[18] ;
    assign n527 = a[18]  & b[18] ;
    assign n528 = ~n526 & ~n527;
    assign n529 = n525 & ~n528;
    assign n530 = ~n525 & n528;
    assign result[18]  = ~n529 & ~n530;
    assign n532 = ~n525 & ~n526;
    assign n533 = ~n527 & ~n532;
    assign n534 = ~a[19]  & ~b[19] ;
    assign n535 = a[19]  & b[19] ;
    assign n536 = ~n534 & ~n535;
    assign n537 = n533 & ~n536;
    assign n538 = ~n533 & n536;
    assign result[19]  = ~n537 & ~n538;
    assign n540 = ~n533 & ~n534;
    assign n541 = ~n535 & ~n540;
    assign n542 = ~a[20]  & ~b[20] ;
    assign n543 = a[20]  & b[20] ;
    assign n544 = ~n542 & ~n543;
    assign n545 = n541 & ~n544;
    assign n546 = ~n541 & n544;
    assign result[20]  = ~n545 & ~n546;
    assign n548 = ~n541 & ~n542;
    assign n549 = ~n543 & ~n548;
    assign n550 = ~a[21]  & ~b[21] ;
    assign n551 = a[21]  & b[21] ;
    assign n552 = ~n550 & ~n551;
    assign n553 = n549 & ~n552;
    assign n554 = ~n549 & n552;
    assign result[21]  = ~n553 & ~n554;
    assign n556 = ~n549 & ~n550;
    assign n557 = ~n551 & ~n556;
    assign n558 = ~a[22]  & ~b[22] ;
    assign n559 = a[22]  & b[22] ;
    assign n560 = ~n558 & ~n559;
    assign n561 = n557 & ~n560;
    assign n562 = ~n557 & n560;
    assign result[22]  = ~n561 & ~n562;
    assign n564 = ~n557 & ~n558;
    assign n565 = ~n559 & ~n564;
    assign n566 = ~a[23]  & ~b[23] ;
    assign n567 = a[23]  & b[23] ;
    assign n568 = ~n566 & ~n567;
    assign n569 = n565 & ~n568;
    assign n570 = ~n565 & n568;
    assign result[23]  = ~n569 & ~n570;
    assign n572 = ~n565 & ~n566;
    assign n573 = ~n567 & ~n572;
    assign n574 = ~a[24]  & ~b[24] ;
    assign n575 = a[24]  & b[24] ;
    assign n576 = ~n574 & ~n575;
    assign n577 = n573 & ~n576;
    assign n578 = ~n573 & n576;
    assign result[24]  = ~n577 & ~n578;
    assign n580 = ~n573 & ~n574;
    assign n581 = ~n575 & ~n580;
    assign n582 = ~a[25]  & ~b[25] ;
    assign n583 = a[25]  & b[25] ;
    assign n584 = ~n582 & ~n583;
    assign n585 = n581 & ~n584;
    assign n586 = ~n581 & n584;
    assign result[25]  = ~n585 & ~n586;
    assign n588 = ~n581 & ~n582;
    assign n589 = ~n583 & ~n588;
    assign n590 = ~a[26]  & ~b[26] ;
    assign n591 = a[26]  & b[26] ;
    assign n592 = ~n590 & ~n591;
    assign n593 = n589 & ~n592;
    assign n594 = ~n589 & n592;
    assign result[26]  = ~n593 & ~n594;
    assign n596 = ~n589 & ~n590;
    assign n597 = ~n591 & ~n596;
    assign n598 = ~a[27]  & ~b[27] ;
    assign n599 = a[27]  & b[27] ;
    assign n600 = ~n598 & ~n599;
    assign n601 = n597 & ~n600;
    assign n602 = ~n597 & n600;
    assign result[27]  = ~n601 & ~n602;
    assign n604 = ~n597 & ~n598;
    assign n605 = ~n599 & ~n604;
    assign n606 = ~a[28]  & ~b[28] ;
    assign n607 = a[28]  & b[28] ;
    assign n608 = ~n606 & ~n607;
    assign n609 = n605 & ~n608;
    assign n610 = ~n605 & n608;
    assign result[28]  = ~n609 & ~n610;
    assign n612 = ~n605 & ~n606;
    assign n613 = ~n607 & ~n612;
    assign n614 = ~a[29]  & ~b[29] ;
    assign n615 = a[29]  & b[29] ;
    assign n616 = ~n614 & ~n615;
    assign n617 = n613 & ~n616;
    assign n618 = ~n613 & n616;
    assign result[29]  = ~n617 & ~n618;
    assign n620 = ~n613 & ~n614;
    assign n621 = ~n615 & ~n620;
    assign n622 = ~a[30]  & ~b[30] ;
    assign n623 = a[30]  & b[30] ;
    assign n624 = ~n622 & ~n623;
    assign n625 = n621 & ~n624;
    assign n626 = ~n621 & n624;
    assign result[30]  = ~n625 & ~n626;
    assign n628 = ~n621 & ~n622;
    assign n629 = ~n623 & ~n628;
    assign n630 = ~a[31]  & ~b[31] ;
    assign n631 = a[31]  & b[31] ;
    assign n632 = ~n630 & ~n631;
    assign n633 = n629 & ~n632;
    assign n634 = ~n629 & n632;
    assign result[31]  = ~n633 & ~n634;
  endmodule

