// int32 add
// deyuan, 09/25/2024

module add_int32(input [31:0] a, input [31:0] b, output [31:0] result);
    assign result = a + b;
endmodule

