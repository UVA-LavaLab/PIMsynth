// 16-bit Signed Integer Min
// Dependencies: gt_int_nbit.v subtractor_1bit_cmp.v, mux_nbit.v
// deyuan, 03/30/2025

module min_int16 #(
    parameter WIDTH = 16,
    parameter IMPL_TYPE = 1
)(
    input [WIDTH-1:0] A,
    input [WIDTH-1:0] B,
    output [WIDTH-1:0] Y,
);

    wire gt;
    gt_int_nbit #(
        .WIDTH(WIDTH),
        .IMPL_TYPE(IMPL_TYPE)
    ) u_gt_int_nbit (
        .A(A),
        .B(B),
        .Y(gt)
    );

    mux_nbit #(.WIDTH(WIDTH)) max_sel ( .A(B), .B(A), .sel(gt), .Y(Y));

endmodule
